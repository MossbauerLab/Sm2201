module dig_machine_ip3601();

endmodule
